module invertebrate (
    input clk,
    input [2:0] reg_1,
    input [2:0] reg_2,
    input [2:0] reg_select,
    input [3:0] alu_op,
    output reg [15:0] alu_result
);
    
endmodule